module odometer_full(AC_STRESS_CLK, SCANOUT_DIN, SCANIN_DIN, SCANIN_CLK, SCANOUT_CLK, RESETB, LOAD, MEAS_TRIG, AC_STRESS_CLK_INT, SCANIN_CLK_INT, SCANOUT_CLK_INT, RESETB_INT, LOAD_INT, MEAS_TRIG_INT, SCANOUT_DOUT, SCANIN_DOUT,VDD,VSS);

	input AC_STRESS_CLK, SCANOUT_DIN, SCANIN_DIN, SCANIN_CLK, SCANOUT_CLK, RESETB, LOAD, MEAS_TRIG,VDD,VSS;
	output AC_STRESS_CLK_INT, SCANIN_CLK_INT, SCANOUT_CLK_INT, RESETB_INT, LOAD_INT, MEAS_TRIG_INT, SCANOUT_DOUT, SCANIN_DOUT;
	
	wire SEL_INV, SEL_NAND, SEL_NOR;
	wire START;
	wire AC_DC,VCO_OUT;
	wire MEAS_STRESS, EN_ROSC, EN_POWR_ROSC_STRESS;
	wire ROSC_STRESS_OUT, ROSC_REF_OUT;

        odometer_meas_ctrl odometer_meas_ctrl(.VCO_OUT(VCO_OUT),.ROSC_STRESS(ROSC_STRESS_OUT), .ROSC_REF(ROSC_REF_OUT), .SEL_INV(SEL_INV), .SEL_NAND(SEL_NAND), .SEL_NOR(SEL_NOR), .START(START), .AC_DC(AC_DC), .VCO(AC_STRESS_CLK), .SCANCHAIN_IN(SCANOUT_DIN), .SCAN_IN(SCANIN_DIN), .SCAN_CLK1(SCANIN_CLK), .SCAN_CLK2(SCANOUT_CLK), .RESETB(RESETB), .LOAD(LOAD), .MEAS_TRIG(MEAS_TRIG), .VCO_INT(AC_STRESS_CLK_INT), .SCAN_CLK1_INT(SCANIN_CLK_INT), .SCAN_CLK2_INT(SCANOUT_CLK_INT), .RESETB_INT(RESETB_INT), .LOAD_INT(LOAD_INT), .MEAS_TRIG_INT(MEAS_TRIG_INT), .SCAN_OUT_INT(SCANOUT_DOUT), .SCANIN_CHECK_INT(SCANIN_DOUT), .MEAS_STRESS(MEAS_STRESS), .EN_ROSC(EN_ROSC), .EN_POWER_ROSC_STRESS(EN_POWER_ROSC_STRESS),.VDD(VDD),.VSS(VSS));

	rosc_block_top_pwr_stress rosc_stress(.SEL_INV(SEL_INV), .SEL_NAND(SEL_NAND), .SEL_NOR(SEL_NOR), .START(START), .AC_DC(AC_DC), .VCO(VCO_OUT), .EN_POWER_ROSC(EN_POWER_ROSC_STRESS), .EN_ROSC(EN_ROSC), .MEAS_STRESS(MEAS_STRESS), .OUT(ROSC_STRESS_OUT));
	
	rosc_block_top_pwr_ref rosc_ref(.SEL_INV(SEL_INV), .SEL_NAND(SEL_NAND), .SEL_NOR(SEL_NOR), .START(MEAS_STRESS), .AC_DC(AC_DC), .VCO(VCO_OUT), .EN_POWER_ROSC(MEAS_STRESS), .EN_ROSC(EN_ROSC), .MEAS_STRESS(MEAS_STRESS), .OUT(ROSC_REF_OUT));

endmodule
